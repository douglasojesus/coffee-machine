module muxA (CLK, S0, S1, S2, S3, SR, SP, SN, VL, M, a);

	or (a, S0, S1, S2, S3, SR, SP, SN, VL);

endmodule